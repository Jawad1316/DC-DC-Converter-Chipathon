** sch_path:
*+ /home/shahid/Desktop/EDA/test/DC_DC_Converter_xschem/1-10-22_xschem/DC_DC_Converter_xschem/DC_DC_Converter/current_pump/current_pump_for_symbol_TB.sch
**.subckt current_pump_for_symbol_TB
X1 UP OUT VDD VSS DN current_pump_for_symbol
C1 OUT GND 20n m=1
V11 UP GND pulse(1.8 0 0 0.01ns 0.01ns 3n 9ns 0)
V3 DN GND pulse(0 1.8 6n 0.01ns 0.01ns 3n 9ns 0)
V1 VDD GND 1.8
V2 VSS GND 0
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/shahid/OSPDKs/sky130A/libs.tech/ngspice/sky130.lib.spice tt




.control
tran 0.1n 50n
plot i(V2) i(V1)
plot v(up) v(dn)

*print @m.xm1.msky130_fd_pr__nfet_01v8
.endc


**** end user architecture code
**.ends

* expanding   symbol:  DC_DC_Converter/current_pump/current_pump_for_symbol.sym # of pins=5
** sym_path:
*+ /home/shahid/Desktop/EDA/test/DC_DC_Converter_xschem/1-10-22_xschem/DC_DC_Converter_xschem/DC_DC_Converter/current_pump/current_pump_for_symbol.sym
** sch_path:
*+ /home/shahid/Desktop/EDA/test/DC_DC_Converter_xschem/1-10-22_xschem/DC_DC_Converter_xschem/DC_DC_Converter/current_pump/current_pump_for_symbol.sch
.subckt current_pump_for_symbol  UP VOUT VDD VSS DN
*.iopin VDD
*.iopin UP
*.iopin DN
*.iopin VSS
*.iopin VOUT
XM1 VOUT DN net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=20 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 VOUT UP net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=60 nf=20 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
R1 net2 VDD sky130_fd_pr__res_generic_m1 W=0.14 L=14.23 m=1
R2 VSS net1 sky130_fd_pr__res_generic_m1 W=0.14 L=11.21 m=1
.ends

.GLOBAL GND
.end
