** sch_path: /home/shahid/Desktop/EDA/test/xschem/Delay_block/Inverter_TB.sch
**.subckt Inverter_TB
X1 VOUT VIN net1 GND inverter
V3 net1 GND 1.8
V5 VIN GND pulse(0 1.8 0 10p 10p 5u 10u 0)
C1 VOUT GND 1p m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/shahid/OSPDKs/sky130A/libs.tech/ngspice/sky130.lib.spice tt




.control
tran 0.5u 50u
plot v(VIN)
plot v(VOUT)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/shahid/Desktop/EDA/test/xschem/inverter.sym
** sch_path: /home/shahid/Desktop/EDA/test/xschem/inverter.sch
.subckt inverter  VOUT VIN VDD VSS
*.iopin VDD
*.iopin VOUT
*.iopin VSS
*.iopin VIN
XM1 VOUT VIN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 VOUT VIN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=12 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
