** sch_path:
*+ /home/shahid/Desktop/EDA/test/1-10-22_xschem/DC_DC_Converter_xschem/DC_DC_Converter/Delay_block_revised/delay_block_stage1_wo_cap.sch
**.subckt delay_block_stage1_wo_cap VDD VSS VIN VOUT
*.iopin VDD
*.iopin VSS
*.iopin VIN
*.iopin VOUT
X_OR1 VDD VSS 1 b net17 OR
X_OR2 VDD VSS 3 d net18 OR
X_OR3 VDD VSS 5 f net19 OR
X_OR4 VDD VSS 7 h net20 OR
X_OR5 VDD VSS net17 net18 ph1 OR
X_OR6 VDD VSS net19 net20 net21 OR
X_OR7 VDD VSS ph1 net21 vin2 OR
X_OR8 VDD VSS VIN vin2 VOUT OR
X13 c net7 VDD VSS Inverter0
X10 net7 net8 VDD VSS Inverter0
X11 4 d VDD VSS Inverter0
X7 b net5 VDD VSS Inverter0
X8 net5 net6 VDD VSS Inverter0
X9 3 c VDD VSS Inverter0
X4 a net3 VDD VSS Inverter0
X5 net3 net4 VDD VSS Inverter0
X6 2 b VDD VSS Inverter0
X1 VIN net1 VDD VSS Inverter0
X2 net1 net2 VDD VSS Inverter0
X3 1 a VDD VSS Inverter0
X12 d net9 VDD VSS Inverter0
X14 net9 net10 VDD VSS Inverter0
X15 5 e VDD VSS Inverter0
X16 e net11 VDD VSS Inverter0
X17 net11 net12 VDD VSS Inverter0
X18 6 f VDD VSS Inverter0
X19 f net13 VDD VSS Inverter0
X20 net13 net14 VDD VSS Inverter0
X21 7 g VDD VSS Inverter0
X22 g net15 VDD VSS Inverter0
X23 net15 net16 VDD VSS Inverter0
X24 8 h VDD VSS Inverter0
X25 net2 1 VDD VSS Inverter0
X26 net4 2 VDD VSS Inverter0
X27 net6 3 VDD VSS Inverter0
X28 net8 4 VDD VSS Inverter0
X29 net10 5 VDD VSS Inverter0
X30 net12 6 VDD VSS Inverter0
X31 net14 7 VDD VSS Inverter0
X32 net16 8 VDD VSS Inverter0
**.ends

* expanding   symbol:  DC_DC_Converter/Delay_block_revised/OR_GATE/OR.sym # of pins=5
** sym_path:
*+ /home/shahid/Desktop/EDA/test/1-10-22_xschem/DC_DC_Converter_xschem/DC_DC_Converter/Delay_block_revised/OR_GATE/OR.sym
** sch_path:
*+ /home/shahid/Desktop/EDA/test/1-10-22_xschem/DC_DC_Converter_xschem/DC_DC_Converter/Delay_block_revised/OR_GATE/OR.sch
.subckt OR  VDD VSS A B OUT
*.iopin VDD
*.iopin VSS
*.iopin A
*.iopin B
*.iopin OUT
XM2 net1 A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM1 net1 B net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM4 net1 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 OUT net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 OUT net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
.ends


* expanding   symbol:  DC_DC_Converter/Delay_block_revised/Inverter_0/Inverter0.sym # of pins=4
** sym_path:
*+ /home/shahid/Desktop/EDA/test/1-10-22_xschem/DC_DC_Converter_xschem/DC_DC_Converter/Delay_block_revised/Inverter_0/Inverter0.sym
** sch_path:
*+ /home/shahid/Desktop/EDA/test/1-10-22_xschem/DC_DC_Converter_xschem/DC_DC_Converter/Delay_block_revised/Inverter_0/Inverter0.sch
.subckt Inverter0  VIN VOUT VDD VSS
*.ipin VIN
*.iopin VDD
*.iopin VSS
*.opin VOUT
XM1 VOUT VIN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 VOUT VIN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
