** sch_path:
*+ /home/shahid/Desktop/EDA/test/DC_DC_Converter_xschem/1-10-22_xschem/DC_DC_Converter_xschem/DC_DC_Converter/Delay_block_revised/AND_GATE/AND_PEX_TB.sch
**.subckt AND_PEX_TB
V2 VDD GND 1.8
V5 VSS GND 0
V1 B GND 1.8
V3 A GND pulse (0 1.8 0 1n 1n 4n 10n 0)
xAND1 VDD VSS A B OUT AND_PEX
**** begin user architecture code


.include ./AND_flatten.spice
.control
tran 0.2n 50n
plot v(OUT) v(A) v(B)
.endc


** manual skywater pdks install (with patches applied)
* .lib /home/shahid/OSPDKs/sky130A/libs.tech/ngspice/models/sky130.lib.spice tt

** opencircuitdesign pdks install
.lib /home/shahid/OSPDKs/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/shahid/OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
