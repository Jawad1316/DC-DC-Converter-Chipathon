** sch_path:
*+ /home/shahid/Desktop/EDA/test/1-10-22_xschem/DC_DC_Converter_xschem/OTHERS/DC_DC_Converter_V7/Non_Overlap_Clk/Non_over_clk_V3.sch
**.subckt Non_over_clk_V3 VDD VSS CLK PH1 PH2
*.iopin VDD
*.iopin VSS
*.iopin CLK
*.iopin PH1
*.iopin PH2
x3 CLK PH1 VSS VSS VDD VDD net3 sky130_fd_sc_hd__nor2_1
x4 net1 VB1 VSS VSS VDD VDD net2 sky130_fd_sc_hd__nor2_1
x6 CLK VSS VSS VDD VDD net1 sky130_fd_sc_hd__clkinv_1
x2 net2 VSS VSS VDD VDD PH1 sky130_fd_sc_hd__clkdlybuf4s50_1
x5 net3 VSS VSS VDD VDD VB1 sky130_fd_sc_hd__clkdlybuf4s50_1
X1 VB1 PH2 VDD VSS Inverter0
**.ends

* expanding   symbol:  DC_DC_Converter/Inverter_0/Inverter0.sym # of pins=4
** sym_path:
*+ /home/shahid/Desktop/EDA/test/1-10-22_xschem/DC_DC_Converter_xschem/DC_DC_Converter/Inverter_0/Inverter0.sym
** sch_path:
*+ /home/shahid/Desktop/EDA/test/1-10-22_xschem/DC_DC_Converter_xschem/DC_DC_Converter/Inverter_0/Inverter0.sch
.subckt Inverter0  VIN VOUT VDD VSS
*.ipin VIN
*.iopin VDD
*.iopin VSS
*.opin VOUT
XM1 VOUT VIN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 VOUT VIN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
