* NGSPICE file created from TopA_flatten.ext - technology: sky130A

.subckt Top_1_PEX VDD VSS SAWTOOTH VREF IBIAS1 OUT1 IBIAS2 IL
X0 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.21275e+15p pd=7.5117e+09u as=1.52741e+15p ps=9.75482e+09u w=1.5e+07u l=150000u
X1 a_5681_22118# a_2807_1109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.56858e+14p ps=2.33496e+09u w=420000u l=150000u
X2 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X3 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X4 VSS a_11826_17500# a_10949_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+13p ps=4.1218e+08u w=8e+06u l=900000u
X5 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X6 a_10711_10879# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=6.96e+12p pd=6.54e+07u as=0p ps=0u w=800000u l=900000u
X7 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.64e+14p ps=1.6528e+09u w=1e+07u l=150000u
X8 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X9 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X10 a_4931_4248# a_2831_3719# a_4511_4248# VDD sky130_fd_pr__pfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X11 VDD a_1901_18557# a_2189_6712# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+13p ps=2.458e+08u w=1.2e+07u l=150000u
X12 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X13 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X14 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X15 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X16 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X17 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X18 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X19 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X20 a_10769_10791# OUT1 VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.59e+07u
X21 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X22 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X23 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X24 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X25 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X26 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X27 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X28 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X29 a_10711_10879# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X30 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X31 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X32 VDD a_5703_18547# a_5991_6702# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+13p ps=2.458e+08u w=1.2e+07u l=150000u
X33 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X34 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X35 a_2435_1206# a_2093_2981# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=3.16e+06u as=0p ps=0u w=500000u l=150000u
X36 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X37 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X38 a_4091_3729# a_2831_3719# a_3671_3729# VSS sky130_fd_pr__nfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X39 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X40 VSS a_12692_11507# a_14220_10933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+12p ps=1.308e+07u w=800000u l=900000u
X41 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X42 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X43 a_11508_10872# VREF a_10949_10879# VSS sky130_fd_pr__nfet_01v8 ad=2.32e+13p pd=1.6464e+08u as=0p ps=0u w=1e+07u l=900000u
X44 a_7907_1338# a_7051_1266# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=150000u
X45 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X46 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X47 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X48 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X49 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X50 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X51 a_2189_6712# a_1901_18557# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.16e+13p pd=8.58e+07u as=0p ps=0u w=4e+06u l=150000u
X52 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X53 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X54 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X55 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X56 a_12750_12001# a_13334_16745# a_13334_16745# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+12p pd=2.116e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=900000u
X57 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X58 a_12692_11507# a_12750_12001# a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=3.48e+12p pd=3.27e+07u as=6.96e+12p ps=6.54e+07u w=800000u l=900000u
X59 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X60 VDD IBIAS1 a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X61 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X62 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X63 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X64 a_6631_1785# a_4957_1270# a_6211_1785# VSS sky130_fd_pr__nfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X65 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X66 a_11508_10872# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X67 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X68 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X69 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X70 a_11508_10872# a_12750_12001# a_12692_11507# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X71 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X72 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X73 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X74 a_9712_6291# a_12750_12001# a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=3.48e+12p pd=3.27e+07u as=0p ps=0u w=800000u l=900000u
X75 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X76 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X77 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X78 VDD IBIAS1 a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X79 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X80 a_11826_17500# a_11814_14752# a_11814_14752# VSS sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.748e+07u as=1.392e+12p ps=1.308e+07u w=800000u l=900000u
X81 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X82 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X83 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X84 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X85 a_11508_10872# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X86 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X87 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X88 a_11508_10872# a_12750_12001# a_12692_11507# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X89 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X90 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X91 a_2189_6712# a_1901_18557# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X92 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X93 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X94 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X95 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X96 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X97 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X98 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X99 VDD IBIAS1 a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X100 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X101 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X102 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X103 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X104 a_11508_10872# VREF a_10949_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X105 a_5791_1785# a_4957_1270# a_5371_1785# VSS sky130_fd_pr__nfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X106 a_10711_10879# a_12750_12001# a_9712_6291# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X107 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X108 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X109 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X110 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X111 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X112 a_10711_10879# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X113 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X114 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X115 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X116 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X117 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X118 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X119 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X120 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X121 a_7021_4248# a_5351_3729# a_6601_4248# VDD sky130_fd_pr__pfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X122 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X123 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X124 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X125 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X126 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X127 a_4117_1789# a_2435_1755# a_3697_1789# VSS sky130_fd_pr__nfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X128 a_7051_1266# a_4957_1270# a_6631_1266# VDD sky130_fd_pr__pfet_01v8 ad=1.247e+11p pd=1.44e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X129 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X130 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X131 a_5761_3729# a_5351_3729# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.494e+11p pd=2.88e+06u as=0p ps=0u w=430000u l=150000u
X132 a_11814_14752# a_11814_14752# a_11826_17500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X133 a_2831_3719# a_3203_3631# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=3.16e+06u as=0p ps=0u w=500000u l=150000u
X134 a_5991_6702# a_5703_18547# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.16e+13p pd=8.58e+07u as=0p ps=0u w=4e+06u l=150000u
X135 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X136 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X137 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X138 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X139 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X140 IBIAS1 IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.658e+07u as=0p ps=0u w=8e+06u l=900000u
X141 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X142 VDD a_5703_18547# a_5991_6702# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X143 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X144 VDD a_1901_18557# a_2189_6712# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X145 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X146 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X147 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X148 a_10711_10879# a_12750_12001# a_9712_6291# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X149 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X150 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X151 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X152 VDD IBIAS1 a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X153 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X154 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X155 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X156 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X157 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X158 a_11508_10872# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X159 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X160 a_1901_18557# a_1839_22225# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+12p pd=2.458e+07u as=0p ps=0u w=1.2e+07u l=150000u
X161 a_11508_10872# VREF a_10949_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X162 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X163 a_8560_7818# a_8560_7818# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X164 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X165 a_1195_24344# a_3203_3631# VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=150000u
X166 a_11508_10872# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X167 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X168 a_6211_1266# a_4957_1270# a_5791_1266# VDD sky130_fd_pr__pfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X169 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X170 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X171 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X172 a_9712_6291# a_12750_12001# a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X173 VDD IBIAS1 a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X174 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X175 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X176 a_17339_1632# a_26051_1314# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X177 a_9712_6291# a_12750_12001# a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X178 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X179 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X180 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X181 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X182 a_9712_6291# a_11814_14752# a_14220_10933# VSS sky130_fd_pr__nfet_01v8 ad=6.96e+11p pd=6.54e+06u as=0p ps=0u w=800000u l=900000u
X183 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X184 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X185 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X186 VDD a_5703_18547# a_5991_6702# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X187 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X188 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X189 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X190 a_11508_10872# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X191 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X192 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X193 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X194 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X195 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X196 a_9712_6291# a_12750_12001# a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X197 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X198 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X199 VDD IBIAS1 a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X200 a_12692_11507# a_12750_12001# a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X201 VDD IBIAS1 a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X202 VDD IBIAS1 a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X203 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X204 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X205 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X206 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X207 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X208 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X209 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X210 VDD a_1901_18557# a_2189_6712# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X211 a_10711_10879# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X212 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X213 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X214 a_10711_10879# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X215 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X216 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X217 VDD a_1901_18557# a_2189_6712# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X218 a_2435_1755# a_2807_1109# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=3.16e+06u as=0p ps=0u w=500000u l=150000u
X219 a_2189_6712# a_1901_18557# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X220 a_12692_11507# a_12750_12001# a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X221 VDD IBIAS1 a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X222 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X223 a_8788_6571# a_8560_7818# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X224 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X225 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X226 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X227 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X228 a_8339_3147# a_7441_3729# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=150000u
X229 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X230 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X231 a_10711_10879# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X232 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X233 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X234 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X235 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X236 a_12692_11507# a_12750_12001# a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X237 VDD a_5681_22118# a_5641_22215# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X238 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X239 a_1901_18557# a_1839_22225# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=150000u
X240 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X241 VSS a_12692_11507# a_14220_10933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X242 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X243 a_3671_3729# a_2831_3719# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X244 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X245 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X246 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X247 VDD a_8618_7721# a_8560_7818# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=500000u
X248 a_6181_4248# a_5351_3729# a_5761_4248# VDD sky130_fd_pr__pfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X249 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X250 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X251 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X252 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X253 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
D0 VSS a_1195_24344# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X254 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X255 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X256 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X257 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X258 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X259 a_12692_11507# a_12750_12001# a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X260 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X261 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X262 a_12692_11507# a_12750_12001# a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X263 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X264 a_7441_3729# a_5351_3729# a_7021_3729# VSS sky130_fd_pr__nfet_01v8 ad=1.247e+11p pd=1.44e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X265 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X266 a_2189_6712# a_1901_18557# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X267 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X268 a_17339_2268# a_26051_2586# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X269 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X270 a_11508_10872# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X271 a_5991_6702# a_5703_18547# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X272 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X273 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X274 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X275 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X276 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X277 a_5703_18547# a_5641_22215# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=150000u
X278 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X279 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X280 a_10711_10879# a_12750_12001# a_9712_6291# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X281 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X282 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X283 a_4537_1789# a_2435_1755# a_4117_1789# VSS sky130_fd_pr__nfet_01v8 ad=2.494e+11p pd=2.88e+06u as=0p ps=0u w=430000u l=150000u
X284 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X285 a_9712_6291# a_11814_14752# a_14220_10933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X286 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X287 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X288 VSS a_12692_11507# a_12688_10937# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+12p ps=1.308e+07u w=800000u l=900000u
X289 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X290 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X291 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X292 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X293 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X294 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X295 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X296 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X297 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X298 a_9712_6291# a_12750_12001# a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X299 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X300 VDD IBIAS1 a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X301 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X302 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X303 VDD IBIAS1 a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X304 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X305 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X306 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X307 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X308 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X309 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X310 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X311 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X312 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X313 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X314 a_6601_3729# a_5351_3729# a_6181_3729# VSS sky130_fd_pr__nfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X315 a_4957_1270# a_2435_1755# a_4537_1270# VDD sky130_fd_pr__pfet_01v8 ad=1.247e+11p pd=1.44e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X316 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X317 a_10711_10879# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X318 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X319 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X320 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X321 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X322 a_12688_10937# a_11814_14752# a_12692_11507# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.96e+11p ps=6.54e+06u w=800000u l=900000u
X323 a_20816_4573# a_9712_6291# VSS sky130_fd_pr__res_xhigh_po_0p35 l=1.819e+07u
X324 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X325 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X326 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X327 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X328 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X329 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X330 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X331 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X332 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X333 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X334 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X335 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X336 a_3697_1789# a_2435_1755# a_3277_1789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X337 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X338 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X339 a_6631_1266# a_4957_1270# a_6211_1266# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X340 a_10711_10879# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X341 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X342 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X343 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X344 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X345 a_2831_3719# a_2141_3069# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X346 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X347 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X348 a_9584_7719# a_8618_7721# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.316e+07u as=0p ps=0u w=3e+06u l=500000u
X349 VSS a_12692_11507# a_14220_10933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X350 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X351 a_9712_6291# a_12750_12001# a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X352 a_10711_10879# a_12750_12001# a_9712_6291# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X353 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X354 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X355 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X356 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X357 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X358 a_11508_10872# a_12750_12001# a_12692_11507# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X359 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X360 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X361 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X362 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X363 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X364 a_4091_4248# a_2831_3719# a_3671_4248# VDD sky130_fd_pr__pfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X365 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X366 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X367 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X368 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X369 VSS a_11826_17500# a_11826_17500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=900000u
X370 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X371 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X372 a_2141_3069# a_2093_2981# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=150000u
X373 VDD a_1901_18557# a_2189_6712# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X374 a_2807_1109# a_8339_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=150000u
X375 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X376 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X377 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X378 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X379 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X380 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X381 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X382 a_10711_10879# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X383 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X384 a_5351_3729# a_2831_3719# a_4931_3729# VSS sky130_fd_pr__nfet_01v8 ad=1.247e+11p pd=1.44e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X385 a_10769_10791# a_26051_1314# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X386 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X387 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X388 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X389 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X390 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X391 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X392 a_5791_1266# a_4957_1270# a_5371_1266# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X393 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X394 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X395 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X396 a_19340_4577# OUT1 VSS sky130_fd_pr__res_xhigh_po_0p35 l=1.47e+06u
X397 a_11814_14752# a_11814_14752# a_11826_17500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X398 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X399 a_3203_3631# a_7907_1338# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=150000u
X400 VSS a_12692_11507# a_12688_10937# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X401 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X402 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X403 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X404 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X405 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X406 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X407 a_10711_10879# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X408 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X409 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X410 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X411 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X412 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X413 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X414 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X415 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X416 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X417 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X418 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X419 a_1879_22128# a_1195_24344# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X420 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X421 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X422 a_17339_3540# a_26051_3222# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X423 a_12692_11507# a_12750_12001# a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X424 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X425 a_7907_1338# a_7051_1266# VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=150000u
X426 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X427 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X428 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X429 a_9712_6291# a_12750_12001# a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X430 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X431 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X432 VDD a_1879_22128# a_1839_22225# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X433 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X434 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X435 a_2435_1755# a_2807_1109# a_2435_1206# VDD sky130_fd_pr__pfet_01v8 ad=1.45e+11p pd=1.58e+06u as=0p ps=0u w=500000u l=150000u
X436 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X437 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X438 a_4511_3729# a_2831_3719# a_4091_3729# VSS sky130_fd_pr__nfet_01v8 ad=2.494e+11p pd=2.88e+06u as=0p ps=0u w=430000u l=150000u
X439 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X440 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X441 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X442 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X443 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X444 IBIAS2 SAWTOOTH a_8618_7721# VSS sky130_fd_pr__nfet_01v8_lvt ad=2.9e+12p pd=2.116e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=700000u
X445 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X446 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X447 a_12692_11507# a_12750_12001# a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X448 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X449 a_5991_6702# a_5703_18547# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X450 VDD a_9584_7719# a_8788_6571# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=500000u
X451 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X452 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X453 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X454 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X455 a_1195_24344# a_3203_3631# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=150000u
X456 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X457 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X458 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X459 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X460 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X461 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X462 a_11826_17500# a_11814_14752# a_11814_14752# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X463 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X464 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X465 a_5681_22118# a_2807_1109# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X466 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X467 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X468 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X469 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X470 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X471 a_11508_10872# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X472 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X473 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X474 a_5761_4248# a_5351_3729# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X475 a_11508_10872# a_12750_12001# a_12692_11507# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X476 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X477 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X478 a_17339_2268# a_26051_1950# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X479 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X480 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X481 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X482 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X483 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X484 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X485 a_10711_10879# a_12750_12001# a_9712_6291# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X486 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X487 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X488 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X489 a_11508_10872# VREF a_10949_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X490 a_10711_10879# a_12750_12001# a_9712_6291# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X491 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X492 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X493 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X494 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X495 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X496 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X497 a_14220_10933# a_11814_14752# a_9712_6291# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X498 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X499 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X500 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X501 VDD a_5703_18547# a_5991_6702# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X502 a_3277_1270# a_2435_1755# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.494e+11p pd=2.88e+06u as=0p ps=0u w=430000u l=150000u
X503 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X504 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X505 a_11508_10872# VREF a_10949_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X506 VSS a_11826_17500# a_10949_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=900000u
X507 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X508 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X509 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X510 a_11508_10872# a_12750_12001# a_12692_11507# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X511 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X512 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X513 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X514 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X515 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X516 a_2141_3069# a_2093_2981# VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=150000u
X517 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X518 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X519 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X520 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X521 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X522 a_5991_6702# a_5703_18547# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X523 a_11508_10872# VREF a_10949_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X524 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X525 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X526 a_11814_14752# a_11814_14752# a_11826_17500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X527 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X528 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X529 VDD IBIAS1 a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X530 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X531 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X532 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X533 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X534 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X535 VSS a_12692_11507# a_12688_10937# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X536 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X537 a_9712_6291# a_12750_12001# a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X538 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X539 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X540 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X541 a_11508_10872# a_12750_12001# a_12692_11507# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X542 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X543 a_5991_6702# a_5703_18547# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X544 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X545 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X546 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X547 a_12688_10937# a_11814_14752# a_12692_11507# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X548 a_10949_10879# a_10769_10791# a_10711_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.32e+13p ps=1.6464e+08u w=1e+07u l=900000u
X549 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X550 a_2831_3719# a_3203_3631# a_2831_4268# VDD sky130_fd_pr__pfet_01v8 ad=1.45e+11p pd=1.58e+06u as=2.9e+11p ps=3.16e+06u w=500000u l=150000u
X551 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X552 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X553 a_2093_2981# a_8788_6571# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X554 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
D1 VSS a_2807_1109# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X555 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X556 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X557 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X558 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X559 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X560 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X561 a_9712_6291# a_12750_12001# a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X562 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X563 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X564 a_10949_10879# a_10769_10791# a_10711_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X565 a_9712_6291# a_10769_10791# sky130_fd_pr__cap_mim_m3_1 l=2.25e+07u w=2.2e+07u
X566 a_5991_6702# a_5703_18547# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X567 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X568 a_11814_14752# a_11814_14752# a_11826_17500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X569 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X570 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X571 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X572 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X573 VDD a_5703_18547# a_5991_6702# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X574 a_11508_10872# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X575 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X576 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X577 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X578 a_10949_10879# a_10769_10791# a_10711_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X579 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X580 a_5991_6702# a_5703_18547# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X581 VDD IBIAS1 a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X582 a_12692_11507# a_12750_12001# a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X583 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X584 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X585 a_3671_4248# a_2831_3719# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X586 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X587 a_2189_6712# a_1901_18557# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X588 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X589 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X590 a_9584_7719# a_9712_6291# IBIAS2 VSS sky130_fd_pr__nfet_01v8_lvt ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=700000u
X591 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X592 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X593 VSS a_1879_22128# a_1839_22225# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X594 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X595 a_10711_10879# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X596 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X597 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X598 a_8339_3147# a_7441_3729# VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=150000u
X599 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X600 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X601 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X602 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X603 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X604 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X605 a_4931_3729# a_2831_3719# a_4511_3729# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X606 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X607 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X608 a_7441_3729# a_5351_3729# a_7021_4248# VDD sky130_fd_pr__pfet_01v8 ad=1.247e+11p pd=1.44e+06u as=0p ps=0u w=430000u l=150000u
X609 VDD IBIAS1 a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X610 a_12692_11507# a_12750_12001# a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X611 VDD IBIAS1 a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X612 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X613 a_2093_2981# a_8788_6571# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=7.25e+11p pd=5.58e+06u as=0p ps=0u w=2.5e+06u l=500000u
X614 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X615 VDD a_1901_18557# a_2189_6712# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X616 a_10711_10879# a_12750_12001# a_9712_6291# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X617 VDD a_5703_18547# a_5991_6702# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X618 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X619 a_10711_10879# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X620 a_11508_10872# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X621 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X622 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X623 a_11508_10872# a_12750_12001# a_12692_11507# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X624 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X625 a_17339_2904# a_26051_3222# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X626 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X627 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X628 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X629 a_11826_17500# a_11814_14752# a_11814_14752# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X630 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X631 a_11826_17500# a_11814_14752# a_11814_14752# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X632 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X633 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X634 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X635 VDD a_9584_7719# a_8618_7721# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.316e+07u w=3e+06u l=500000u
X636 a_9712_6291# a_12750_12001# a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X637 a_20816_4573# a_10769_10791# sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=3.4e+06u
X638 VDD IBIAS1 a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X639 VSS a_5681_22118# a_5641_22215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X640 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X641 VDD IBIAS1 a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X642 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X643 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X644 a_12692_11507# a_11814_14752# a_12688_10937# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X645 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X646 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X647 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X648 a_5371_1785# a_4957_1270# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X649 VDD a_13334_16745# VSS sky130_fd_pr__res_high_po_0p35 l=1e+06u
X650 a_1879_22128# a_1195_24344# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X651 a_11508_10872# a_12750_12001# a_12692_11507# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X652 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X653 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X654 a_12692_11507# a_12750_12001# a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X655 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X656 VDD a_5703_18547# a_5991_6702# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X657 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X658 VDD IBIAS1 a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X659 VDD a_1901_18557# a_2189_6712# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X660 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X661 a_6601_4248# a_5351_3729# a_6181_4248# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X662 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X663 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X664 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X665 a_11814_14752# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.658e+07u as=0p ps=0u w=8e+06u l=900000u
X666 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X667 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X668 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X669 a_14220_10933# a_12692_11507# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X670 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X671 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X672 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X673 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X674 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X675 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X676 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X677 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X678 a_2189_6712# a_1901_18557# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X679 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X680 a_10949_10879# a_10769_10791# a_10711_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X681 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X682 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X683 VDD a_1901_18557# a_2189_6712# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X684 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X685 a_4117_1270# a_2435_1755# a_3697_1270# VDD sky130_fd_pr__pfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X686 a_9712_6291# a_12750_12001# a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X687 VDD IBIAS1 a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X688 a_10949_10879# a_10769_10791# a_10711_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X689 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X690 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X691 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X692 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X693 VDD IBIAS1 a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X694 a_9584_7719# a_9584_7719# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X695 a_4957_1270# a_2435_1755# a_4537_1789# VSS sky130_fd_pr__nfet_01v8 ad=1.247e+11p pd=1.44e+06u as=0p ps=0u w=430000u l=150000u
X696 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X697 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X698 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X699 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X700 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X701 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X702 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X703 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X704 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X705 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X706 a_10711_10879# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X707 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X708 VSS a_11826_17500# a_10949_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=900000u
X709 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X710 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X711 a_12688_10937# a_12692_11507# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X712 a_14220_10933# a_11814_14752# a_9712_6291# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X713 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X714 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X715 VSS a_26051_3858# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X716 a_10711_10879# a_12750_12001# a_9712_6291# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X717 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X718 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X719 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X720 VDD IBIAS1 a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X721 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X722 a_2189_6712# a_1901_18557# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X723 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X724 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X725 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X726 a_7021_3729# a_5351_3729# a_6601_3729# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X727 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X728 a_5351_3729# a_2831_3719# a_4931_4248# VDD sky130_fd_pr__pfet_01v8 ad=1.247e+11p pd=1.44e+06u as=0p ps=0u w=430000u l=150000u
X729 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X730 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X731 a_10711_10879# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X732 a_11508_10872# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X733 VDD a_5703_18547# a_5991_6702# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X734 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X735 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X736 VDD IBIAS1 a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X737 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X738 a_9712_6291# a_12750_12001# a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X739 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X740 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X741 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X742 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X743 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X744 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X745 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X746 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X747 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X748 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X749 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X750 VSS a_11826_17500# a_10949_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=900000u
X751 a_2807_1109# a_8339_3147# VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=150000u
X752 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X753 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X754 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X755 a_12692_11507# a_11814_14752# a_12688_10937# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X756 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X757 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X758 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X759 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X760 a_10949_10879# a_10769_10791# a_10711_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X761 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X762 VDD a_5703_18547# a_5991_6702# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X763 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X764 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X765 VDD IBIAS1 a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X766 a_2189_6712# a_1901_18557# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X767 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X768 a_2435_1755# a_2093_2981# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X769 VDD IBIAS1 a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X770 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X771 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X772 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X773 a_2831_4268# a_2141_3069# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X774 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X775 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X776 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X777 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X778 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X779 a_14220_10933# a_12692_11507# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X780 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X781 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X782 a_4511_4248# a_2831_3719# a_4091_4248# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X783 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X784 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X785 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X786 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X787 a_7051_1266# a_4957_1270# a_6631_1785# VSS sky130_fd_pr__nfet_01v8 ad=1.247e+11p pd=1.44e+06u as=0p ps=0u w=430000u l=150000u
X788 a_17339_2904# a_26051_2586# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X789 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X790 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X791 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X792 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X793 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X794 a_3203_3631# a_7907_1338# VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=150000u
X795 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X796 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X797 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X798 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X799 a_8618_7721# a_8618_7721# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X800 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X801 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X802 a_13334_16745# VSS VSS sky130_fd_pr__res_high_po_0p35 l=1e+06u
X803 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X804 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X805 VDD IBIAS1 a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X806 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X807 a_12692_11507# a_12750_12001# a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X808 a_12692_11507# a_12750_12001# a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X809 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X810 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X811 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X812 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X813 VDD a_1901_18557# a_2189_6712# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X814 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X815 a_9712_6291# a_12750_12001# a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X816 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X817 a_12750_12001# a_12750_12001# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=900000u
X818 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X819 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X820 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X821 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X822 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X823 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X824 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X825 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X826 a_12688_10937# a_12692_11507# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X827 a_14220_10933# a_11814_14752# a_9712_6291# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X828 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X829 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X830 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X831 a_10949_10879# a_10769_10791# a_10711_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X832 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X833 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X834 a_12692_11507# a_12750_12001# a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X835 a_12692_11507# a_12750_12001# a_11508_10872# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X836 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X837 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X838 a_6211_1785# a_4957_1270# a_5791_1785# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X839 a_5991_6702# a_5703_18547# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X840 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X841 a_10711_10879# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X842 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X843 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X844 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X845 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X846 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X847 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X848 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X849 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X850 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X851 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X852 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X853 a_10711_10879# a_12750_12001# a_9712_6291# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X854 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X855 a_11508_10872# VREF a_10949_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X856 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X857 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X858 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X859 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X860 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X861 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X862 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X863 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X864 a_6181_3729# a_5351_3729# a_5761_3729# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X865 a_4537_1270# a_2435_1755# a_4117_1270# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X866 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X867 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X868 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X869 a_2189_6712# a_1901_18557# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X870 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X871 a_19340_4577# a_10769_10791# sky130_fd_pr__cap_mim_m3_1 l=9.8e+06u w=9.9e+06u
X872 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X873 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X874 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X875 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X876 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X877 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X878 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X879 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X880 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X881 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X882 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X883 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X884 a_17339_3540# a_26051_3858# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X885 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X886 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X887 a_5991_6702# a_5703_18547# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X888 a_3277_1789# a_2435_1755# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X889 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X890 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X891 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X892 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X893 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X894 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X895 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X896 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X897 a_10949_10879# a_10769_10791# a_10711_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X898 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X899 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X900 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X901 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X902 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X903 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X904 a_5991_6702# a_5703_18547# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X905 VSS a_11826_17500# a_10949_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=900000u
X906 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X907 a_11826_17500# a_11814_14752# a_11814_14752# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X908 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X909 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X910 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X911 a_11508_10872# a_12750_12001# a_12692_11507# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X912 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X913 a_2189_6712# a_1901_18557# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X914 VDD a_5703_18547# a_5991_6702# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X915 a_3697_1270# a_2435_1755# a_3277_1270# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X916 a_11814_14752# a_11814_14752# a_11826_17500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X917 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X918 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X919 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X920 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X921 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X922 a_11508_10872# VREF a_10949_10879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X923 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X924 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X925 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X926 a_17339_1632# a_26051_1950# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X927 a_10711_10879# a_12750_12001# a_9712_6291# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X928 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X929 VDD a_1901_18557# a_2189_6712# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X930 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X931 a_9712_6291# a_12750_12001# a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X932 a_9712_6291# a_12750_12001# a_10711_10879# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X933 IL a_5991_6702# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X934 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X935 a_11508_10872# a_12750_12001# a_12692_11507# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X936 VSS a_5991_6702# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X937 a_5703_18547# a_5641_22215# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+12p pd=2.458e+07u as=0p ps=0u w=1.2e+07u l=150000u
X938 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X939 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X940 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X941 a_12688_10937# a_11814_14752# a_12692_11507# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X942 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X943 VDD a_2189_6712# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X944 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X945 a_5371_1266# a_4957_1270# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X946 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X947 IL a_2189_6712# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
.ends

