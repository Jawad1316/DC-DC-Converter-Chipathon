* NGSPICE file created from Top.ext - technology: sky130A

.subckt Top_PEX VDD VSS VREF IL VH IBIAS1 VL IBIAS2 ENABLE BIAS3 OUT BIAS4 SAWTOOTH
X0 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=1.64874e+15p pd=1.0707e+10u as=1.21275e+15p ps=7.5117e+09u w=1.5e+07u l=150000u
X1 a_71263_34662# a_70433_34133# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.98891e+14p ps=2.7043e+09u w=420000u l=150000u
X2 VSS a_71263_34662# a_72241_31805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.84e+06u w=420000u l=150000u
X3 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X4 a_10308_7770# a_8208_7760# a_9888_7770# VSS sky130_fd_pr__nfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X5 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X6 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X7 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.64e+14p ps=1.6528e+09u w=1e+07u l=150000u
X8 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X9 VDD IBIAS1 a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.96e+12p ps=6.54e+07u w=800000u l=900000u
X10 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X11 VDD a_11080_22588# a_11368_10743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+13p ps=2.458e+08u w=1.2e+07u l=150000u
X12 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X13 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X14 BIAS3 VH a_56243_36303# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+12p pd=2.116e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X15 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X16 a_68185_14789# a_68093_13516# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X17 a_18065_14978# a_17191_18793# a_18069_15548# VSS sky130_fd_pr__nfet_01v8 ad=1.392e+12p pd=1.308e+07u as=6.96e+11p ps=6.54e+06u w=800000u l=900000u
X18 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X19 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X20 a_18065_14978# a_18069_15548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X21 a_82606_36983# a_82288_8250# OUT VDD sky130_fd_pr__pfet_01v8 ad=1.077e+13p pd=7.318e+07u as=9.9e+12p ps=6.66e+07u w=3e+06u l=150000u
X22 OUT a_82654_36220# a_82702_36308# VSS sky130_fd_pr__nfet_01v8 ad=3.59e+12p pd=2.918e+07u as=3.3e+12p ps=2.66e+07u w=1e+06u l=150000u
X23 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X24 a_70383_18394# a_67084_14777# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.392e+12p pd=1.424e+07u as=0p ps=0u w=600000u l=150000u
X25 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X26 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X27 VDD a_7278_22598# a_7566_10753# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+13p ps=2.458e+08u w=1.2e+07u l=150000u
X28 VSS a_17203_21541# a_16326_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+13p ps=4.1218e+08u w=8e+06u l=900000u
X29 VDD ENABLE a_55365_29869# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.96e+11p ps=7.12e+06u w=600000u l=150000u
X30 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X31 OUT a_82288_8250# a_82606_36983# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X32 a_82702_36308# a_82654_36220# OUT VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_11368_10743# a_11080_22588# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.16e+13p pd=8.58e+07u as=0p ps=0u w=4e+06u l=150000u
X34 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X35 a_85910_23842# a_73171_11284# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X36 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X37 a_73881_31122# a_73071_32334# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.392e+12p pd=1.424e+07u as=0p ps=0u w=600000u l=150000u
X38 a_73811_14325# a_73007_13942# a_73821_14854# VDD sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=7.12e+06u as=1.392e+12p ps=1.424e+07u w=600000u l=150000u
X39 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X40 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X41 VSS a_58085_30619# a_57725_29899# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.872e+11p ps=5.68e+06u w=420000u l=150000u
X42 a_69386_13417# a_69018_11991# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X43 a_67446_13401# a_67084_14777# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
R0 a_82702_36308# VSS sky130_fd_pr__res_generic_m1 w=140000u l=1.121e+07u
X44 a_73007_13942# a_72177_14863# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X45 a_66305_31041# a_56275_30688# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X46 a_26193_8614# a_15089_10332# VSS sky130_fd_pr__res_xhigh_po_0p35 l=1.819e+07u
X47 VDD a_82000_20095# a_82288_8250# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+13p ps=2.458e+08u w=1.2e+07u l=150000u
X48 a_72187_13230# a_71183_13646# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.392e+12p pd=1.424e+07u as=0p ps=0u w=600000u l=150000u
X49 a_16326_14920# a_16146_14832# a_16088_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.32e+13p ps=1.6464e+08u w=1e+07u l=900000u
X50 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X51 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X52 a_16885_14913# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X53 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X54 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X55 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X56 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X57 a_70369_17191# a_66125_10752# a_70379_15558# VDD sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=7.12e+06u as=1.392e+12p ps=1.424e+07u w=600000u l=150000u
X58 a_73071_32334# a_72241_31805# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X59 a_15089_10332# a_18127_16042# a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=3.48e+12p pd=3.27e+07u as=6.96e+12p ps=6.54e+07u w=800000u l=900000u
X60 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X61 a_67066_26921# VSS sky130_fd_pr__cap_mim_m3_2 l=1.4e+07u w=1.4e+07u
X62 a_73821_14854# a_73011_16066# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X63 VDD a_11080_22588# a_11368_10743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X64 a_67056_12029# a_66217_12025# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X65 a_18069_15548# a_18127_16042# a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=3.48e+12p pd=3.27e+07u as=0p ps=0u w=800000u l=900000u
X66 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X67 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X68 VDD a_66225_26923# a_66185_27020# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X69 a_67084_14777# a_66245_14773# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X70 a_82702_36308# a_82654_36220# OUT VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X71 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X72 VDD a_56185_37833# a_58223_37543# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.25e+11p ps=5.58e+06u w=2.5e+06u l=1e+06u
X73 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X74 a_16088_14920# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X75 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X76 a_9468_8289# a_8208_7760# a_9048_8289# VDD sky130_fd_pr__pfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X77 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X78 a_70433_34133# a_66213_29768# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.84e+06u as=0p ps=0u w=420000u l=150000u
D0 VSS a_81183_36165# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X79 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X80 VSS a_17203_21541# a_16326_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=900000u
X81 a_7470_7022# a_14165_10612# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X82 VSS a_11058_26159# a_11018_26256# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X83 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X84 a_10308_8289# a_8208_7760# a_9888_8289# VDD sky130_fd_pr__pfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X85 a_15089_10332# a_18127_16042# a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X86 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X87 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X88 VDD IBIAS1 a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X89 a_18069_15548# a_18127_16042# a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X90 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X91 VDD a_68127_10617# a_68087_10714# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X92 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X93 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X94 a_70363_13646# a_68127_10617# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.392e+12p pd=1.424e+07u as=0p ps=0u w=600000u l=150000u
X95 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X96 VDD a_11080_22588# a_11368_10743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X97 a_24717_8618# OUT VSS sky130_fd_pr__res_xhigh_po_0p35 l=1.47e+06u
X98 VDD a_66125_10752# a_68968_10615# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X99 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X100 a_16088_14920# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X101 a_16088_14920# a_18127_16042# a_15089_10332# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X102 a_16088_14920# a_18127_16042# a_15089_10332# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X103 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X104 a_70443_34662# a_67144_31045# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.392e+12p pd=1.424e+07u as=0p ps=0u w=600000u l=150000u
X105 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X106 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X107 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X108 a_82288_8250# a_82000_20095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.16e+13p pd=8.58e+07u as=0p ps=0u w=4e+06u l=150000u
X109 OUT a_82654_36220# a_82702_36308# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X110 a_16885_14913# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X111 a_16088_14920# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X112 a_16088_14920# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X113 a_22716_5673# a_31428_5355# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X114 a_66217_12025# a_66153_13500# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X115 a_16885_14913# a_18127_16042# a_18069_15548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X116 a_16885_14913# VREF a_16326_14920# VSS sky130_fd_pr__nfet_01v8 ad=2.32e+13p pd=1.6464e+08u as=0p ps=0u w=1e+07u l=900000u
X117 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X118 a_70413_29385# a_69446_29685# a_70423_29914# VDD sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=7.12e+06u as=1.392e+12p ps=1.424e+07u w=600000u l=150000u
X119 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X120 VSS a_66185_27020# a_69028_26883# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X121 a_14961_11760# a_13995_11762# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.316e+07u as=0p ps=0u w=3e+06u l=500000u
X122 VSS a_18069_15548# a_18065_14978# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X123 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X124 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X125 a_69446_29685# a_69078_28259# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X126 a_72411_27552# a_56275_30688# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.392e+12p pd=1.424e+07u as=0p ps=0u w=600000u l=150000u
X127 a_15089_10332# a_18127_16042# a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X128 VDD IBIAS1 a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X129 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X130 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X131 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X132 a_85932_20271# a_85870_23939# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=150000u
X133 a_72241_31805# a_71259_32538# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X134 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X135 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X136 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X137 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X138 VSS a_66225_26923# a_66185_27020# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X139 a_13937_11859# a_13937_11859# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X140 a_73881_31122# a_73071_32334# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X141 a_70409_28711# a_69506_31063# a_70419_27078# VDD sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=7.12e+06u as=1.392e+12p ps=1.424e+07u w=600000u l=150000u
X142 a_16088_14920# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X143 a_16088_14920# a_18127_16042# a_15089_10332# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X144 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X145 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X146 a_73231_27552# a_72401_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X147 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X148 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X149 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X150 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X151 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X152 a_67116_28297# a_66277_28293# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X153 a_16885_14913# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X154 a_16885_14913# a_18127_16042# a_18069_15548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X155 a_57207_36187# OUT BIAS3 VSS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=1e+06u
X156 a_70433_34133# a_66213_29768# a_70443_34662# VDD sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=7.12e+06u as=0p ps=0u w=600000u l=150000u
X157 a_11978_7770# a_10728_7770# a_11558_7770# VSS sky130_fd_pr__nfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X158 a_72191_16066# a_71203_18394# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.392e+12p pd=1.424e+07u as=0p ps=0u w=600000u l=150000u
X159 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X160 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X161 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X162 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X163 a_9494_5830# a_7812_5796# a_9074_5830# VSS sky130_fd_pr__nfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X164 VDD a_85932_20271# a_82654_36220# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+13p ps=2.458e+08u w=1.2e+07u l=150000u
X165 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X166 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X167 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X168 VSS a_73071_32334# a_73871_30593# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.84e+06u w=420000u l=150000u
X169 a_15089_10332# a_18127_16042# a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X170 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X171 a_11588_5826# a_10334_5311# a_11168_5826# VSS sky130_fd_pr__nfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X172 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X173 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X174 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X175 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X176 VDD IBIAS1 a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X177 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X178 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X179 a_70383_18394# a_67084_14777# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X180 IBIAS1 IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.658e+07u as=0p ps=0u w=8e+06u l=900000u
X181 a_82654_36220# a_85932_20271# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.16e+13p pd=8.58e+07u as=0p ps=0u w=4e+06u l=150000u
X182 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X183 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X184 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X185 a_70349_12443# a_69446_14795# a_70359_10810# VDD sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=7.12e+06u as=1.392e+12p ps=1.424e+07u w=600000u l=150000u
X186 a_11368_10743# a_11080_22588# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X187 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X188 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X189 OUT a_82654_36220# a_82702_36308# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X190 a_7566_10753# a_7278_22598# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.16e+13p pd=8.58e+07u as=0p ps=0u w=4e+06u l=150000u
X191 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X192 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X193 a_72247_29498# a_71243_29914# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.392e+12p pd=1.424e+07u as=0p ps=0u w=600000u l=150000u
X194 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X195 VDD a_82000_20095# a_82288_8250# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X196 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X197 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X198 a_17191_18793# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.658e+07u as=0p ps=0u w=8e+06u l=900000u
X199 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X200 a_68179_11987# VSS sky130_fd_pr__cap_mim_m3_2 l=1.4e+07u w=1.4e+07u
X201 a_82288_8250# a_82000_20095# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X202 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X203 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X204 a_72353_26935# a_73871_30593# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X205 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X206 a_69446_14795# a_69024_14793# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X207 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X208 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X209 a_73821_14854# a_73011_16066# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X210 a_70383_18394# a_67084_14777# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X211 a_66245_14773# a_58547_30718# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X212 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X213 VDD a_7278_22598# a_7566_10753# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X214 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X215 a_16885_14913# a_18127_16042# a_18069_15548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X216 a_70373_17865# a_66153_13500# a_70383_18394# VDD sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=7.12e+06u as=0p ps=0u w=600000u l=150000u
X217 a_71259_32538# a_70429_33459# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X218 a_70353_13117# a_69386_13417# a_70363_13646# VDD sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=7.12e+06u as=0p ps=0u w=600000u l=150000u
X219 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X220 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X221 a_22716_6309# a_31428_5991# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X222 a_70359_10810# a_68133_13419# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X223 a_72293_10667# a_73811_14325# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X224 VDD IBIAS1 a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X225 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X226 a_72237_31131# a_71239_27790# a_72247_29498# VDD sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=7.12e+06u as=0p ps=0u w=600000u l=150000u
X227 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X228 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X229 a_72351_11284# a_58547_30718# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.392e+12p pd=1.424e+07u as=0p ps=0u w=600000u l=150000u
X230 a_19597_14974# a_18069_15548# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.392e+12p pd=1.308e+07u as=0p ps=0u w=800000u l=900000u
D1 VSS a_6572_28385# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X231 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X232 a_72251_32334# a_71263_34662# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.392e+12p pd=1.424e+07u as=0p ps=0u w=600000u l=150000u
X233 a_10334_5311# a_7812_5796# a_9914_5311# VDD sky130_fd_pr__pfet_01v8 ad=1.247e+11p pd=1.44e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X234 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X235 a_73871_30593# a_73067_30210# a_73881_31122# VDD sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=7.12e+06u as=0p ps=0u w=600000u l=150000u
X236 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X237 a_11978_8289# a_10728_7770# a_11558_8289# VDD sky130_fd_pr__pfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X238 a_69446_14795# a_69024_14793# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X239 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X240 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X241 a_11368_10743# a_11080_22588# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X242 a_17203_21541# a_17191_18793# a_17191_18793# VSS sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.748e+07u as=1.392e+12p ps=1.308e+07u w=800000u l=900000u
X243 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X244 a_72241_31805# a_71259_32538# a_72251_32334# VDD sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=7.12e+06u as=0p ps=0u w=600000u l=150000u
X245 a_68245_31057# a_68153_29784# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X246 VDD a_66253_29671# a_66213_29768# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X247 a_15089_10332# a_18127_16042# a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X248 a_7566_10753# a_7278_22598# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X249 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X250 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X251 VDD a_67418_10653# a_67006_10653# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X252 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X253 VDD IBIAS1 a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X254 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X255 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X256 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X257 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X258 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X259 VDD a_7278_22598# a_7566_10753# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X260 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X261 a_82654_36220# a_85932_20271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X262 VDD a_11080_22588# a_11368_10743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X263 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X264 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X265 a_16088_14920# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X266 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X267 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X268 VSS a_67478_26921# a_67066_26921# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X269 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X270 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X271 a_72241_31805# a_71259_32538# a_72251_32334# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X272 a_16885_14913# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X273 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X274 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X275 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X276 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X277 a_7812_5247# a_7470_7022# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=3.16e+06u as=0p ps=0u w=500000u l=150000u
X278 a_82654_36220# a_85932_20271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X279 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X280 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X281 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X282 a_70443_34662# a_67144_31045# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X283 a_70379_15558# a_67056_12029# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X284 a_57725_29899# ENABLE a_57637_29899# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.84e+06u w=420000u l=150000u
X285 a_70433_34133# a_66213_29768# a_70443_34662# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X286 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X287 a_72191_16066# a_71203_18394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X288 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X289 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X290 VSS a_67506_29669# a_67094_29669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X291 a_8654_5311# a_7812_5796# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.494e+11p pd=2.88e+06u as=0p ps=0u w=430000u l=150000u
X292 VDD a_68133_13419# a_68093_13516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X293 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X294 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X295 a_11058_26159# a_8184_5150# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X296 VDD a_7278_22598# a_7566_10753# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X297 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X298 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X299 a_67144_31045# a_66305_31041# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X300 a_16088_14920# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X301 a_71199_16270# a_70369_17191# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X302 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X303 VSS a_67084_14777# a_70373_17865# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.84e+06u w=420000u l=150000u
X304 a_7256_26169# a_6572_28385# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X305 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X306 a_70419_27078# a_68193_29687# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X307 a_10748_5307# a_10334_5311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.494e+11p pd=2.88e+06u as=0p ps=0u w=430000u l=150000u
X308 VSS a_68127_10617# a_70353_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.84e+06u w=420000u l=150000u
X309 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X310 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X311 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X312 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X313 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X314 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X315 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X316 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X317 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X318 VDD IBIAS1 a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X319 VSS a_18069_15548# a_18065_14978# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X320 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X321 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X322 VDD a_11058_26159# a_11018_26256# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X323 a_71239_27790# a_70409_28711# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X324 a_13716_7188# a_12818_7770# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=150000u
X325 VDD a_7256_26169# a_7216_26266# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X326 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X327 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X328 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X329 a_72181_15537# a_71199_16270# a_72191_16066# VDD sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=7.12e+06u as=0p ps=0u w=600000u l=150000u
X330 a_18065_14978# a_17191_18793# a_18069_15548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X331 a_73067_30210# a_72237_31131# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X332 a_66277_28293# a_66213_29768# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X333 a_72187_13230# a_71183_13646# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X334 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X335 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X336 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X337 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X338 VSS a_55813_30589# a_55453_29869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.872e+11p ps=5.68e+06u w=420000u l=150000u
X339 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X340 VSS a_67006_10653# a_66165_10655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X341 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X342 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X343 a_11138_7770# a_10728_7770# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.494e+11p pd=2.88e+06u as=0p ps=0u w=430000u l=150000u
X344 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X345 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X346 a_55813_30589# a_58169_33911# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X347 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X348 a_8208_7760# a_8580_7672# a_8208_8309# VDD sky130_fd_pr__pfet_01v8 ad=1.45e+11p pd=1.58e+06u as=2.9e+11p ps=3.16e+06u w=500000u l=150000u
X349 a_71183_13646# a_70353_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X350 a_71203_18394# a_70373_17865# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X351 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X352 VDD ENABLE a_57637_29899# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.96e+11p ps=7.12e+06u w=600000u l=150000u
X353 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X354 a_66277_28293# a_66213_29768# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X355 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X356 a_70439_31826# a_67116_28297# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.392e+12p pd=1.424e+07u as=0p ps=0u w=600000u l=150000u
X357 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X358 a_72353_26935# a_73871_30593# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X359 a_72177_14863# a_71179_11522# a_72187_13230# VDD sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=7.12e+06u as=0p ps=0u w=600000u l=150000u
X360 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X361 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X362 a_18065_14978# a_17191_18793# a_18069_15548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X363 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X364 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X365 a_72351_11284# a_58547_30718# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X366 a_15089_10332# a_18127_16042# a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X367 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X368 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X369 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X370 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X371 a_18069_15548# a_18127_16042# a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X372 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X373 a_58547_30718# a_57637_29899# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X374 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X375 a_11368_10743# a_11080_22588# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X376 a_71259_32538# a_70429_33459# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X377 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X378 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X379 a_7566_10753# a_7278_22598# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X380 a_70379_15558# a_67056_12029# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X381 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X382 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X383 a_16146_14832# OUT VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.59e+07u
X384 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X385 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X386 a_70349_12443# a_69446_14795# a_70359_10810# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X387 a_68179_11987# a_68087_10714# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X388 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X389 a_55453_29869# ENABLE a_55365_29869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.84e+06u w=420000u l=150000u
X390 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X391 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X392 a_13995_11762# a_13995_11762# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.316e+07u as=0p ps=0u w=3e+06u l=500000u
X393 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X394 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X395 VSS a_56179_37031# a_56179_37031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X396 VSS a_69028_26883# a_68187_26885# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X397 VDD IBIAS1 a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X398 a_15089_10332# a_18127_16042# a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X399 VDD a_82000_20095# a_82288_8250# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X400 a_18127_16042# a_18127_16042# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+12p pd=2.116e+07u as=0p ps=0u w=5e+06u l=900000u
X401 a_72341_10755# a_72293_10667# a_72351_11284# VDD sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=7.12e+06u as=0p ps=0u w=600000u l=150000u
X402 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X403 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X404 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X405 a_18069_15548# a_18127_16042# a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X406 OUT a_82288_8250# a_82606_36983# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X407 a_72241_31805# a_71259_32538# a_72251_32334# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X408 a_70413_29385# a_69446_29685# a_70423_29914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X409 a_16146_14832# a_31428_5355# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X410 a_18069_15548# a_18127_16042# a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X411 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X412 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X413 a_17203_21541# a_17191_18793# a_17191_18793# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X414 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X415 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X416 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X417 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X418 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X419 a_11368_10743# a_11080_22588# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X420 a_73871_30593# a_73067_30210# a_73881_31122# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X421 a_12818_7770# a_10728_7770# a_12398_7770# VSS sky130_fd_pr__nfet_01v8 ad=1.247e+11p pd=1.44e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X422 VSS a_71203_18394# a_72181_15537# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.84e+06u w=420000u l=150000u
X423 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X424 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X425 VSS a_67066_26921# a_66225_26923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X426 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X427 a_16885_14913# a_18127_16042# a_18069_15548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X428 a_7566_10753# a_7278_22598# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X429 VSS a_68193_29687# a_68153_29784# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X430 a_11138_8289# a_10728_7770# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.494e+11p pd=2.88e+06u as=0p ps=0u w=430000u l=150000u
X431 a_70373_17865# a_66153_13500# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X432 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X433 a_12428_5307# a_10334_5311# a_12008_5826# VSS sky130_fd_pr__nfet_01v8 ad=1.247e+11p pd=1.44e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X434 a_70353_13117# a_69386_13417# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X435 VSS a_17203_21541# a_16326_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=900000u
X436 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X437 VSS a_69446_29685# a_69034_29685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X438 a_68968_10615# VSS sky130_fd_pr__cap_mim_m3_2 l=1.4e+07u w=1.4e+07u
X439 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X440 a_69084_31061# a_68245_31057# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X441 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X442 a_73871_30593# a_73067_30210# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X443 VDD IBIAS1 a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X444 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X445 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X446 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X447 VSS a_7256_26169# a_7216_26266# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X448 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X449 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X450 OUT a_82288_8250# a_82606_36983# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X451 a_57153_35149# VL BIAS4 VSS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=2.9e+12p ps=2.116e+07u w=5e+06u l=1e+06u
X452 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X453 a_82702_36308# a_82654_36220# OUT VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X454 a_18069_15548# a_18127_16042# a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X455 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X456 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X457 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X458 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X459 VSS a_17203_21541# a_16326_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=900000u
X460 a_68245_31057# VSS sky130_fd_pr__cap_mim_m3_2 l=1.4e+07u w=1.4e+07u
X461 VDD a_7278_22598# a_7566_10753# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X462 a_82606_36983# a_82288_8250# OUT VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X463 a_72401_27023# a_72353_26935# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.84e+06u as=0p ps=0u w=420000u l=150000u
X464 a_22716_7581# a_31428_7263# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X465 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X466 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X467 VSS a_71243_29914# a_72237_31131# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.84e+06u w=420000u l=150000u
X468 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X469 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X470 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X471 a_70363_13646# a_68127_10617# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X472 a_16885_14913# a_18127_16042# a_18069_15548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X473 VDD ENABLE a_57637_29899# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X474 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X475 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X476 a_16326_14920# a_16146_14832# a_16088_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X477 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X478 a_70439_31826# a_67116_28297# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X479 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X480 VDD a_82000_20095# a_82288_8250# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X481 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X482 a_69078_28259# a_68239_28255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X483 a_70419_27078# a_68193_29687# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X484 VSS a_18069_15548# a_18065_14978# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X485 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X486 a_58547_30718# a_57637_29899# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X487 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X488 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X489 a_17203_21541# a_17191_18793# a_17191_18793# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X490 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X491 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X492 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X493 a_11368_10743# a_11080_22588# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X494 a_8208_7760# a_8580_7672# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=3.16e+06u as=0p ps=0u w=500000u l=150000u
X495 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X496 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X497 a_70423_29914# a_68187_26885# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X498 a_72411_27552# a_56275_30688# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X499 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X500 VDD a_85932_20271# a_82654_36220# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X501 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X502 a_7566_10753# a_7278_22598# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X503 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X504 VDD a_67446_13401# a_67034_13401# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X505 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X506 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X507 a_16326_14920# a_16146_14832# a_16088_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X508 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X509 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X510 a_70353_13117# a_69386_13417# a_70363_13646# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X511 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X512 VSS a_58085_30619# a_57725_29899# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X513 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X514 VSS a_58547_30718# a_72341_10755# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.84e+06u w=420000u l=150000u
X515 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X516 VSS a_56125_34399# a_56131_33597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X517 a_71243_29914# a_70413_29385# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X518 a_12818_7770# a_10728_7770# a_12398_8289# VDD sky130_fd_pr__pfet_01v8 ad=1.247e+11p pd=1.44e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X519 a_73067_30210# a_72237_31131# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X520 a_19597_14974# a_18069_15548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X521 VDD a_82000_20095# a_82288_8250# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X522 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X523 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X524 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X525 a_7518_7110# a_7470_7022# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=150000u
X526 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X527 OUT a_82288_8250# a_82606_36983# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X528 a_82702_36308# a_82654_36220# OUT VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X529 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X530 a_70413_29385# a_69446_29685# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.84e+06u as=0p ps=0u w=420000u l=150000u
X531 VDD a_13995_11762# a_13937_11859# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=500000u
X532 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X533 a_82606_36983# a_82288_8250# OUT VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X534 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X535 a_13716_7188# a_12818_7770# VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=150000u
X536 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X537 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X538 a_56275_30688# a_55365_29869# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X539 a_73871_30593# a_73067_30210# a_73881_31122# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X540 a_72237_31131# a_71239_27790# a_72247_29498# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X541 a_72401_27023# a_72353_26935# a_72411_27552# VDD sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=7.12e+06u as=0p ps=0u w=600000u l=150000u
X542 a_82654_36220# a_85932_20271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X543 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X544 a_82288_8250# a_82000_20095# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X545 VDD a_67006_10653# a_66165_10655# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X546 a_73811_14325# a_73007_13942# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.84e+06u as=0p ps=0u w=420000u l=150000u
X547 a_67116_28297# a_66277_28293# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X548 a_67034_13401# VSS sky130_fd_pr__cap_mim_m3_2 l=1.4e+07u w=1.4e+07u
X549 VDD a_85932_20271# a_82654_36220# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X550 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X551 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X552 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X553 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X554 VDD a_68968_10615# a_68127_10617# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X555 a_82000_20095# a_81938_23763# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=150000u
X556 VDD a_58085_30619# a_57637_29899# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X557 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X558 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X559 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X560 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X561 a_72181_15537# a_71199_16270# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X562 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X563 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X564 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X565 a_73171_11284# a_72341_10755# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X566 a_15089_10332# a_18127_16042# a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X567 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X568 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X569 a_82606_36983# a_82288_8250# OUT VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X570 OUT a_82654_36220# a_82702_36308# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X571 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X572 a_73821_14854# a_73011_16066# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X573 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X574 VSS a_31428_7899# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X575 a_71179_11522# a_70349_12443# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X576 a_16885_14913# VREF a_16326_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X577 VDD a_82000_20095# a_82288_8250# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X578 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X579 VDD a_66193_13403# a_66153_13500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X580 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X581 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X582 a_9494_5311# a_7812_5796# a_9074_5311# VDD sky130_fd_pr__pfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X583 a_70373_17865# a_66153_13500# a_70383_18394# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X584 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X585 VDD IBIAS1 a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X586 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X587 a_14961_11760# a_15089_10332# IBIAS2 VSS sky130_fd_pr__nfet_01v8_lvt ad=1.45e+12p pd=1.058e+07u as=2.9e+12p ps=2.116e+07u w=5e+06u l=700000u
X588 a_70409_28711# a_69506_31063# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.84e+06u as=0p ps=0u w=420000u l=150000u
X589 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X590 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X591 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X592 a_11588_5307# a_10334_5311# a_11168_5307# VDD sky130_fd_pr__pfet_01v8 ad=2.494e+11p pd=2.88e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X593 a_19597_14974# a_17191_18793# a_15089_10332# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.96e+11p ps=6.54e+06u w=800000u l=900000u
X594 VSS a_67094_29669# a_66253_29671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X595 VDD a_85932_20271# a_82654_36220# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X596 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X597 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X598 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X599 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X600 VDD a_85932_20271# a_82654_36220# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X601 a_9888_7770# a_8208_7760# a_9468_7770# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X602 a_82288_8250# a_82000_20095# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X603 a_72191_16066# a_71203_18394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X604 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X605 VSS a_56125_34399# a_56125_34399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X606 a_72237_31131# a_71239_27790# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X607 a_70413_29385# a_69446_29685# a_70423_29914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X608 a_72177_14863# a_71179_11522# a_72187_13230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X609 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X610 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X611 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X612 a_72411_27552# a_56275_30688# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X613 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X614 a_68185_14789# a_68093_13516# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X615 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X616 OUT a_82654_36220# a_82702_36308# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X617 a_71183_13646# a_70353_13117# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X618 a_71203_18394# a_70373_17865# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X619 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X620 a_16885_14913# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X621 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X622 a_10728_7770# a_8208_7760# a_10308_7770# VSS sky130_fd_pr__nfet_01v8 ad=1.247e+11p pd=1.44e+06u as=0p ps=0u w=430000u l=150000u
X623 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X624 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X625 VDD a_56243_36303# a_56179_37031# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X626 a_69028_26883# VSS sky130_fd_pr__cap_mim_m3_2 l=1.4e+07u w=1.4e+07u
X627 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X628 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X629 VDD IBIAS1 a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X630 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X631 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X632 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X633 a_73231_27552# a_72401_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X634 a_19597_14974# a_17191_18793# a_15089_10332# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X635 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X636 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X637 a_67506_29669# a_67144_31045# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X638 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X639 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X640 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X641 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X642 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X643 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X644 a_73811_14325# a_73007_13942# a_73821_14854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X645 VDD a_7278_22598# a_7566_10753# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X646 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X647 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X648 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X649 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X650 a_82654_36220# a_85932_20271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X651 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X652 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X653 a_81183_36165# a_73231_27552# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X654 a_11368_10743# a_11080_22588# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X655 a_73071_32334# a_72241_31805# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X656 a_18069_15548# a_17191_18793# a_18065_14978# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X657 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X658 a_72341_10755# a_72293_10667# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X659 VSS a_56179_37031# a_56185_37833# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X660 a_11058_26159# a_8184_5150# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X661 a_7566_10753# a_7278_22598# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X662 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X663 a_17191_18793# a_17191_18793# a_17203_21541# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X664 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X665 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X666 a_7518_7110# a_7470_7022# VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=150000u
X667 a_7256_26169# a_6572_28385# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X668 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X669 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X670 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X671 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X672 a_70353_13117# a_69386_13417# a_70363_13646# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X673 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X674 a_73881_31122# a_73071_32334# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X675 a_57207_36187# a_56243_36303# VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.16e+06u as=0p ps=0u w=1.5e+06u l=500000u
X676 a_58169_33911# a_56131_33597# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X677 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X678 a_85910_23842# a_73171_11284# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X679 a_82288_8250# a_82000_20095# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X680 a_67084_14777# a_66245_14773# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X681 VSS a_18069_15548# a_19597_14974# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X682 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X683 VDD a_68187_26885# a_68147_26982# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X684 VSS a_68127_10617# a_68087_10714# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X685 a_70433_34133# a_66213_29768# a_70443_34662# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X686 VDD a_58085_30619# a_57637_29899# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X687 VDD a_66185_27020# a_69028_26883# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X688 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X689 a_70439_31826# a_67116_28297# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X690 a_18069_15548# a_18127_16042# a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X691 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X692 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X693 a_16326_14920# a_16146_14832# a_16088_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X694 OUT a_82654_36220# a_82702_36308# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X695 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X696 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X697 a_72351_11284# a_58547_30718# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X698 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X699 a_72401_27023# a_72353_26935# a_72411_27552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X700 a_9888_8289# a_8208_7760# a_9468_8289# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X701 a_16088_14920# a_18127_16042# a_15089_10332# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X702 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X703 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X704 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X705 a_11080_22588# a_11018_26256# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+12p pd=2.458e+07u as=0p ps=0u w=1.2e+07u l=150000u
X706 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X707 a_16885_14913# a_18127_16042# a_18069_15548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X708 a_71263_34662# a_70433_34133# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X709 VDD a_56189_35133# a_56125_34399# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X710 a_57153_35149# a_56189_35133# VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.16e+06u as=0p ps=0u w=1.5e+06u l=500000u
X711 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X712 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X713 a_10728_7770# a_8208_7760# a_10308_8289# VDD sky130_fd_pr__pfet_01v8 ad=1.247e+11p pd=1.44e+06u as=0p ps=0u w=430000u l=150000u
X714 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X715 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X716 a_68239_28255# a_68147_26982# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X717 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X718 VDD a_82000_20095# a_82288_8250# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X719 a_24717_8618# a_16146_14832# sky130_fd_pr__cap_mim_m3_1 l=9.8e+06u w=9.9e+06u
X720 a_15089_10332# a_18127_16042# a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X721 VDD a_85932_20271# a_82654_36220# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X722 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X723 a_7812_5796# a_8184_5150# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=3.16e+06u as=0p ps=0u w=500000u l=150000u
X724 VSS a_68133_13419# a_70349_12443# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.84e+06u w=420000u l=150000u
X725 VDD IBIAS1 a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X726 a_72181_15537# a_71199_16270# a_72191_16066# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X727 a_66305_31041# a_56275_30688# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X728 a_68974_13417# VSS sky130_fd_pr__cap_mim_m3_2 l=1.4e+07u w=1.4e+07u
X729 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X730 a_6572_28385# a_8580_7672# VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=150000u
X731 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X732 a_66277_28293# VSS sky130_fd_pr__cap_mim_m3_2 l=1.4e+07u w=1.4e+07u
X733 VDD IBIAS1 a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X734 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X735 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X736 a_16088_14920# a_18127_16042# a_15089_10332# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X737 a_82702_36308# a_82654_36220# OUT VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X738 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X739 VSS a_66193_13403# a_66153_13500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X740 a_16885_14913# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X741 a_16885_14913# a_18127_16042# a_18069_15548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X742 a_70373_17865# a_66153_13500# a_70383_18394# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X743 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X744 VDD a_67506_29669# a_67094_29669# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X745 VSS a_73011_16066# a_73811_14325# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X746 VSS a_67446_13401# a_67034_13401# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X747 a_13284_5379# a_12428_5307# VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=150000u
X748 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X749 VSS a_69034_29685# a_68193_29687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X750 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X751 a_70359_10810# a_68133_13419# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X752 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X753 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X754 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X755 a_15089_10332# a_18127_16042# a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X756 VDD IBIAS1 a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X757 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X758 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X759 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X760 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X761 a_72237_31131# a_71239_27790# a_72247_29498# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X762 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X763 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X764 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X765 a_82654_36220# a_85932_20271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X766 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X767 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X768 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X769 a_18065_14978# a_18069_15548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X770 a_16088_14920# a_18127_16042# a_15089_10332# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X771 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X772 a_71179_11522# a_70349_12443# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X773 VDD a_68974_13417# a_68133_13419# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X774 a_70373_17865# a_66153_13500# a_70383_18394# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X775 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X776 a_16088_14920# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X777 a_17191_18793# a_17191_18793# a_17203_21541# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X778 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X779 a_9914_5830# a_7812_5796# a_9494_5830# VSS sky130_fd_pr__nfet_01v8 ad=2.494e+11p pd=2.88e+06u as=0p ps=0u w=430000u l=150000u
X780 VDD a_58169_33911# a_55813_30589# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.25e+11p ps=5.58e+06u w=2.5e+06u l=1e+06u
X781 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X782 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X783 a_69018_11991# a_68179_11987# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X784 a_70379_15558# a_67056_12029# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X785 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X786 a_67006_10653# VSS sky130_fd_pr__cap_mim_m3_2 l=1.4e+07u w=1.4e+07u
X787 VSS a_68968_10615# a_68127_10617# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X788 a_12008_5826# a_10334_5311# a_11588_5826# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X789 VDD a_11080_22588# a_11368_10743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X790 a_69506_31063# a_69084_31061# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X791 VSS a_67056_12029# a_70369_17191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.84e+06u w=420000u l=150000u
X792 a_85932_20271# a_85870_23939# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+12p pd=2.458e+07u as=0p ps=0u w=1.2e+07u l=150000u
X793 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X794 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X795 a_22716_6945# a_31428_7263# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X796 a_70349_12443# a_69446_14795# a_70359_10810# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X797 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X798 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X799 VDD a_11080_22588# a_11368_10743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X800 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X801 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X802 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X803 VDD a_69386_13417# a_68974_13417# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X804 VDD a_58223_37543# a_58085_30619# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.25e+11p ps=5.58e+06u w=2.5e+06u l=1e+06u
X805 a_16088_14920# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X806 a_72341_10755# a_72293_10667# a_72351_11284# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X807 a_16088_14920# a_18127_16042# a_15089_10332# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X808 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X809 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X810 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X811 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X812 a_82702_36308# a_82654_36220# OUT VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X813 a_72241_31805# a_71259_32538# a_72251_32334# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X814 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X815 a_67056_12029# a_66217_12025# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X816 VDD a_67034_13401# a_66193_13403# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X817 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X818 a_72353_26935# a_73871_30593# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X819 a_9048_7770# a_8208_7760# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.494e+11p pd=2.88e+06u as=0p ps=0u w=430000u l=150000u
X820 VSS a_66125_10752# a_68968_10615# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X821 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X822 a_16326_14920# a_16146_14832# a_16088_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X823 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X824 a_70423_29914# a_68187_26885# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X825 a_72247_29498# a_71243_29914# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X826 VDD a_14961_11760# a_14165_10612# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=500000u
X827 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X828 a_11080_22588# a_11018_26256# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=150000u
X829 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X830 a_8580_7672# a_13284_5379# VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=150000u
X831 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X832 a_69018_11991# a_68179_11987# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X833 a_82288_8250# a_82000_20095# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X834 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X835 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X836 a_67418_10653# a_67056_12029# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X837 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X838 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X839 a_82654_36220# a_85932_20271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X840 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X841 VSS a_56275_30688# a_72401_27023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X842 a_73171_11284# a_72341_10755# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X843 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X844 a_73071_32334# a_72241_31805# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X845 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X846 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X847 VSS a_17203_21541# a_16326_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=900000u
X848 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X849 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X850 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X851 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X852 VSS a_55813_30589# a_55453_29869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X853 a_71199_16270# a_70369_17191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X854 BIAS4 OUT a_56189_35133# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X855 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X856 VSS a_71183_13646# a_72177_14863# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.84e+06u w=420000u l=150000u
X857 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X858 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X859 VDD a_81978_23666# a_81938_23763# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X860 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X861 VDD IBIAS1 a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X862 a_70349_12443# a_69446_14795# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X863 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X864 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X865 a_70433_34133# a_66213_29768# a_70443_34662# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X866 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X867 a_16088_14920# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X868 a_70369_17191# a_66125_10752# a_70379_15558# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X869 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X870 a_57725_29899# ENABLE a_57637_29899# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X871 a_58547_30718# a_57637_29899# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X872 VDD a_14961_11760# a_13995_11762# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X873 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X874 a_70439_31826# a_67116_28297# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X875 a_16885_14913# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X876 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X877 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X878 a_15089_10332# a_16146_14832# sky130_fd_pr__cap_mim_m3_1 l=2.25e+07u w=2.2e+07u
X879 a_72181_15537# a_71199_16270# a_72191_16066# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X880 a_70419_27078# a_68193_29687# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X881 a_72187_13230# a_71183_13646# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X882 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X883 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X884 a_70409_28711# a_69506_31063# a_70419_27078# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X885 a_73231_27552# a_72401_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X886 VDD a_82000_20095# a_82288_8250# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X887 a_8184_5150# a_13716_7188# VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=150000u
X888 a_68179_11987# a_68087_10714# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X889 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X890 VDD a_11080_22588# a_11368_10743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X891 VDD a_68193_29687# a_68153_29784# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X892 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X893 a_12428_5307# a_10334_5311# a_12008_5307# VDD sky130_fd_pr__pfet_01v8 ad=1.247e+11p pd=1.44e+06u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X894 VSS a_68133_13419# a_68093_13516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X895 a_16885_14913# VREF a_16326_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X896 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X897 VDD a_55813_30589# a_55365_29869# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X898 a_71239_27790# a_70409_28711# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X899 VDD a_11080_22588# a_11368_10743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X900 VDD a_69446_29685# a_69034_29685# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X901 a_69446_29685# a_69078_28259# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X902 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X903 a_16088_14920# a_18127_16042# a_15089_10332# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X904 VSS a_68187_26885# a_70413_29385# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X905 a_81978_23666# a_81183_36165# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X906 a_16088_14920# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X907 a_66245_14773# a_58547_30718# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X908 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X909 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X910 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X911 a_9048_8289# a_8208_7760# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X912 a_70413_29385# a_69446_29685# a_70423_29914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X913 a_16885_14913# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X914 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X915 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X916 a_73011_16066# a_72181_15537# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=3.56e+06u as=0p ps=0u w=600000u l=150000u
X917 a_15089_10332# a_18127_16042# a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X918 a_15089_10332# a_18127_16042# a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X919 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X920 VSS a_68187_26885# a_68147_26982# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X921 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X922 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X923 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X924 a_17203_21541# a_17191_18793# a_17191_18793# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X925 VDD IBIAS1 a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X926 a_72177_14863# a_71179_11522# a_72187_13230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X927 a_18069_15548# a_18127_16042# a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X928 a_70369_17191# a_66125_10752# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X929 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X930 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X931 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X932 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X933 a_70379_15558# a_67056_12029# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X934 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X935 VDD a_11080_22588# a_11368_10743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X936 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X937 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X938 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X939 a_17203_21541# a_17191_18793# a_17191_18793# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X940 a_16088_14920# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X941 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X942 a_82288_8250# a_82000_20095# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X943 a_55453_29869# ENABLE a_55365_29869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X944 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X945 a_15089_10332# a_17191_18793# a_19597_14974# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X946 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X947 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X948 a_73007_13942# a_72177_14863# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X949 a_15089_10332# a_18127_16042# a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X950 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X951 a_70429_33459# a_66185_27020# a_70439_31826# VDD sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=7.12e+06u as=0p ps=0u w=600000u l=150000u
X952 a_71243_29914# a_70413_29385# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X953 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X954 VSS a_68193_29687# a_70409_28711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X955 a_72341_10755# a_72293_10667# a_72351_11284# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X956 a_73811_14325# a_73007_13942# a_73821_14854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X957 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X958 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X959 a_73067_30210# a_72237_31131# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X960 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X961 VDD IBIAS1 a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X962 a_18069_15548# a_18127_16042# a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X963 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X964 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X965 a_72293_10667# a_73811_14325# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X966 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X967 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X968 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X969 a_16088_14920# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X970 a_14961_11760# a_14961_11760# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X971 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X972 a_16088_14920# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X973 a_66305_31041# VSS sky130_fd_pr__cap_mim_m3_2 l=1.4e+07u w=1.4e+07u
X974 a_70369_17191# a_66125_10752# a_70379_15558# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X975 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X976 a_16885_14913# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X977 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X978 a_67478_26921# a_67116_28297# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X979 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X980 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X981 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X982 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X983 a_11558_7770# a_10728_7770# a_11138_7770# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X984 a_72177_14863# a_71179_11522# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X985 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X986 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X987 a_82606_36983# a_82288_8250# OUT VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X988 VDD a_69028_26883# a_68187_26885# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X989 a_9074_5830# a_7812_5796# a_8654_5830# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X990 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X991 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X992 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X993 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X994 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X995 a_69024_14793# a_68185_14789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X996 a_73011_16066# a_72181_15537# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X997 a_18069_15548# a_17191_18793# a_18065_14978# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X998 a_67144_31045# a_66305_31041# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X999 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1000 a_11168_5826# a_10334_5311# a_10748_5826# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.494e+11p ps=2.88e+06u w=430000u l=150000u
X1001 a_16885_14913# VREF a_16326_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X1002 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1003 a_68239_28255# VSS sky130_fd_pr__cap_mim_m3_2 l=1.4e+07u w=1.4e+07u
X1004 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1005 a_70423_29914# a_68187_26885# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1006 a_14165_10612# a_13937_11859# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X1007 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1008 VDD a_7278_22598# a_7566_10753# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X1009 a_16088_14920# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1010 a_56275_30688# a_55365_29869# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1011 a_71239_27790# a_70409_28711# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X1012 a_70429_33459# a_66185_27020# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.84e+06u as=0p ps=0u w=420000u l=150000u
X1013 VSS a_81978_23666# a_81938_23763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1014 a_69034_29685# VSS sky130_fd_pr__cap_mim_m3_2 l=1.4e+07u w=1.4e+07u
X1015 a_67446_13401# a_67084_14777# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X1016 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1017 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1018 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1019 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1020 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1021 a_18069_15548# a_18127_16042# a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1022 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1023 VDD ENABLE a_55365_29869# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1024 a_70419_27078# a_68193_29687# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1025 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1026 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1027 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1028 VDD a_57207_36187# a_56243_36303# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.16e+06u w=1.5e+06u l=500000u
X1029 VSS a_17203_21541# a_17203_21541# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=900000u
X1030 a_82654_36220# a_85932_20271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1031 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1032 a_70443_34662# a_67144_31045# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1033 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1034 VDD a_56131_33597# a_58169_33911# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.25e+11p ps=5.58e+06u w=2.5e+06u l=1e+06u
X1035 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1036 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1037 a_68239_28255# a_68147_26982# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1038 a_16885_14913# a_18127_16042# a_18069_15548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1039 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1040 a_7812_5796# a_8184_5150# a_7812_5247# VDD sky130_fd_pr__pfet_01v8 ad=1.45e+11p pd=1.58e+06u as=0p ps=0u w=500000u l=150000u
X1041 a_22716_6945# a_31428_6627# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X1042 VDD a_67094_29669# a_66253_29671# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X1043 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1044 VSS a_67034_13401# a_66193_13403# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1045 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1046 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1047 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1048 VDD a_57153_35149# a_56189_35133# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.16e+06u w=1.5e+06u l=500000u
X1049 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1050 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1051 a_18127_16042# a_18711_20786# a_18711_20786# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=900000u
X1052 a_70353_13117# a_69386_13417# a_70363_13646# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1053 a_82606_36983# a_82288_8250# OUT VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1054 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1055 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1056 a_56131_33597# a_57153_35149# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1057 a_70429_33459# a_66185_27020# a_70439_31826# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1058 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1059 a_70359_10810# a_68133_13419# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1060 a_18069_15548# a_18127_16042# a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1061 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1062 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1063 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1064 a_70409_28711# a_69506_31063# a_70419_27078# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1065 a_73007_13942# a_72177_14863# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X1066 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
R1 a_82606_36983# VDD sky130_fd_pr__res_generic_m1 w=140000u l=1.423e+07u
X1067 a_11558_8289# a_10728_7770# a_11138_8289# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X1068 a_7278_22598# a_7216_26266# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+12p pd=2.458e+07u as=0p ps=0u w=1.2e+07u l=150000u
X1069 a_16885_14913# a_18127_16042# a_18069_15548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1070 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1071 a_73871_30593# a_73067_30210# a_73881_31122# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1072 a_72401_27023# a_72353_26935# a_72411_27552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1073 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1074 a_69386_13417# a_69018_11991# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X1075 a_71183_13646# a_70353_13117# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1076 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1077 VDD IBIAS1 a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1078 a_82288_8250# a_82000_20095# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1079 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1080 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1081 VDD a_67478_26921# a_67066_26921# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X1082 VDD a_18711_20786# VSS sky130_fd_pr__res_high_po_0p35 l=1e+06u
X1083 a_82654_36220# a_85932_20271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1084 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1085 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1086 a_82288_8250# a_82000_20095# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1087 a_70383_18394# a_67084_14777# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1088 VDD a_7278_22598# a_7566_10753# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X1089 a_16326_14920# a_16146_14832# a_16088_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X1090 a_70363_13646# a_68127_10617# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1091 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1092 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1093 VDD a_7278_22598# a_7566_10753# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X1094 OUT a_82288_8250# a_82606_36983# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1095 VDD IBIAS1 a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1096 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1097 a_73811_14325# a_73007_13942# a_73821_14854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1098 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1099 a_8184_5150# a_13716_7188# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=150000u
X1100 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1101 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1102 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1103 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1104 a_69506_31063# a_69084_31061# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1105 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1106 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1107 a_72247_29498# a_71243_29914# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1108 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1109 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1110 VDD IBIAS1 a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1111 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1112 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1113 a_68185_14789# VSS sky130_fd_pr__cap_mim_m3_2 l=1.4e+07u w=1.4e+07u
X1114 a_72251_32334# a_71263_34662# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1115 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1116 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1117 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1118 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1119 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1120 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1121 OUT a_82288_8250# a_82606_36983# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1122 a_82702_36308# a_82654_36220# OUT VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1123 VDD a_7278_22598# a_7566_10753# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X1124 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1125 a_7566_10753# a_7278_22598# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1126 a_69084_31061# a_68245_31057# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1127 a_26193_8614# a_16146_14832# sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=3.4e+06u
X1128 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1129 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1130 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1131 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1132 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1133 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1134 VSS a_67418_10653# a_67006_10653# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1135 a_67418_10653# a_67056_12029# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1136 a_71203_18394# a_70373_17865# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1137 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1138 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1139 a_56243_36303# a_56243_36303# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1140 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1141 VDD a_82000_20095# a_82288_8250# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X1142 a_82288_8250# a_82000_20095# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1143 a_11368_10743# a_11080_22588# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1144 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1145 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1146 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1147 a_72251_32334# a_71263_34662# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1148 a_7566_10753# a_7278_22598# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1149 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1150 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1151 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1152 a_16885_14913# VREF a_16326_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X1153 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1154 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1155 OUT a_82288_8250# a_82606_36983# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1156 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
D2 VSS a_8184_5150# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
D3 VSS a_73171_11284# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X1157 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1158 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1159 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1160 VDD a_57153_35149# a_57153_35149# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1161 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1162 a_22716_7581# a_31428_7899# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X1163 a_72181_15537# a_71199_16270# a_72191_16066# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1164 a_70443_34662# a_67144_31045# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1165 a_81978_23666# a_81183_36165# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1166 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1167 a_72401_27023# a_72353_26935# a_72411_27552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1168 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1169 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1170 VDD a_57207_36187# a_57207_36187# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1171 a_7278_22598# a_7216_26266# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=150000u
X1172 VDD a_69034_29685# a_68193_29687# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X1173 a_8208_8309# a_7518_7110# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1174 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1175 a_17191_18793# a_17191_18793# a_17203_21541# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1176 a_17191_18793# a_17191_18793# a_17203_21541# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1177 VSS a_85910_23842# a_85870_23939# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1178 a_16885_14913# VREF a_16326_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X1179 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1180 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1181 a_71179_11522# a_70349_12443# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1182 a_73821_14854# a_73011_16066# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1183 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1184 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1185 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1186 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1187 VDD a_66165_10655# a_66125_10752# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X1188 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1189 OUT a_82288_8250# a_82606_36983# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1190 a_82702_36308# a_82654_36220# OUT VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1191 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1192 a_58085_30619# a_58223_37543# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X1193 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1194 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1195 a_9914_5311# a_7812_5796# a_9494_5311# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X1196 a_72293_10667# a_73811_14325# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1197 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1198 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1199 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1200 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1201 VDD a_85932_20271# a_82654_36220# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X1202 a_11368_10743# a_11080_22588# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1203 a_72191_16066# a_71203_18394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1204 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1205 VDD IBIAS1 a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1206 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1207 a_12008_5307# a_10334_5311# a_11588_5307# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X1208 VDD a_85932_20271# a_82654_36220# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X1209 a_7566_10753# a_7278_22598# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1210 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1211 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1212 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1213 a_6572_28385# a_8580_7672# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=150000u
X1214 a_82654_36220# a_85932_20271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1215 VDD a_85932_20271# a_82654_36220# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X1216 a_69078_28259# a_68239_28255# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1217 a_66217_12025# a_66153_13500# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X1218 a_15089_10332# a_18127_16042# a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1219 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1220 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1221 a_22716_5673# a_31428_5991# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X1222 a_15089_10332# a_17191_18793# a_19597_14974# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1223 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1224 VDD a_82000_20095# a_82288_8250# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X1225 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1226 a_18069_15548# a_18127_16042# a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1227 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1228 a_82606_36983# a_82288_8250# OUT VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1229 OUT a_82654_36220# a_82702_36308# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1230 a_10334_5311# a_7812_5796# a_9914_5830# VSS sky130_fd_pr__nfet_01v8 ad=1.247e+11p pd=1.44e+06u as=0p ps=0u w=430000u l=150000u
X1231 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1232 VSS a_66253_29671# a_66213_29768# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1233 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1234 a_13284_5379# a_12428_5307# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=150000u
X1235 a_72187_13230# a_71183_13646# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1236 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1237 a_70429_33459# a_66185_27020# a_70439_31826# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1238 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1239 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1240 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1241 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1242 a_17191_18793# a_17191_18793# a_17203_21541# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1243 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1244 a_72341_10755# a_72293_10667# a_72351_11284# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1245 a_71263_34662# a_70433_34133# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1246 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1247 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1248 a_12398_7770# a_10728_7770# a_11978_7770# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X1249 a_71199_16270# a_70369_17191# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1250 VDD a_11080_22588# a_11368_10743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X1251 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1252 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1253 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1254 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1255 VDD IBIAS1 a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1256 a_15089_10332# a_18127_16042# a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1257 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1258 a_73881_31122# a_73071_32334# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1259 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1260 a_18069_15548# a_18127_16042# a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1261 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1262 a_82606_36983# a_82288_8250# OUT VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1263 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1264 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1265 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1266 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1267 OUT a_82654_36220# a_82702_36308# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1268 a_66217_12025# VSS sky130_fd_pr__cap_mim_m3_2 l=1.4e+07u w=1.4e+07u
X1269 a_70359_10810# a_68133_13419# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1270 a_18069_15548# a_18127_16042# a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1271 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1272 a_70423_29914# a_68187_26885# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1273 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1274 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1275 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1276 a_82000_20095# a_81938_23763# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+12p pd=2.458e+07u as=0p ps=0u w=1.2e+07u l=150000u
X1277 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1278 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1279 a_72351_11284# a_58547_30718# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1280 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1281 a_72251_32334# a_71263_34662# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1282 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1283 OUT a_82288_8250# a_82606_36983# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1284 a_71243_29914# a_70413_29385# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1285 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1286 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1287 a_16326_14920# a_16146_14832# a_16088_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X1288 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1289 VDD IBIAS1 a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1290 a_8654_5830# a_7812_5796# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X1291 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1292 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1293 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1294 a_18711_20786# VSS VSS sky130_fd_pr__res_high_po_0p35 l=1e+06u
X1295 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1296 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1297 a_70349_12443# a_69446_14795# a_70359_10810# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1298 a_10748_5826# a_10334_5311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X1299 a_18069_15548# a_18127_16042# a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1300 a_58223_37543# a_56185_37833# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X1301 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1302 a_82606_36983# a_82288_8250# OUT VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1303 OUT a_82654_36220# a_82702_36308# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1304 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1305 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1306 a_8580_7672# a_13284_5379# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=150000u
X1307 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1308 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1309 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1310 a_8208_7760# a_7518_7110# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1311 a_16885_14913# a_18127_16042# a_18069_15548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1312 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1313 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1314 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1315 VSS a_18069_15548# a_19597_14974# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1316 VDD a_85932_20271# a_82654_36220# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=150000u
X1317 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1318 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1319 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1320 a_16326_14920# a_16146_14832# a_16088_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X1321 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1322 VDD a_55813_30589# a_55365_29869# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1323 a_66245_14773# VSS sky130_fd_pr__cap_mim_m3_2 l=1.4e+07u w=1.4e+07u
X1324 a_70369_17191# a_66125_10752# a_70379_15558# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1325 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1326 a_22716_6309# a_31428_6627# VSS sky130_fd_pr__res_xhigh_po_0p35 l=4.14e+07u
X1327 VSS a_68974_13417# a_68133_13419# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1328 a_12398_8289# a_10728_7770# a_11978_8289# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X1329 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1330 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1331 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1332 a_82606_36983# a_82288_8250# OUT VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1333 a_73171_11284# a_72341_10755# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1334 a_16088_14920# a_18127_16042# a_15089_10332# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1335 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1336 OUT a_82654_36220# a_82702_36308# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1337 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1338 a_68245_31057# a_68153_29784# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1339 VDD a_85910_23842# a_85870_23939# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X1340 VSS a_67116_28297# a_70429_33459# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1341 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1342 VSS a_18069_15548# a_19597_14974# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1343 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1344 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1345 a_16885_14913# IBIAS1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1346 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1347 a_67478_26921# a_67116_28297# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1348 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1349 VDD a_67066_26921# a_66225_26923# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
X1350 VSS a_69386_13417# a_68974_13417# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1351 a_56189_35133# a_56189_35133# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1352 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1353 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1354 a_56275_30688# a_55365_29869# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X1355 a_72237_31131# a_71239_27790# a_72247_29498# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1356 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1357 a_19597_14974# a_17191_18793# a_15089_10332# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1358 a_16885_14913# VREF a_16326_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X1359 VSS a_67144_31045# a_70433_34133# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1360 a_67506_29669# a_67144_31045# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1361 a_56185_37833# a_57207_36187# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1362 a_69024_14793# a_68185_14789# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1363 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1364 a_16088_14920# a_18127_16042# a_15089_10332# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1365 a_70363_13646# a_68127_10617# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1366 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1367 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1368 OUT a_82288_8250# a_82606_36983# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1369 a_82702_36308# a_82654_36220# OUT VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1370 IBIAS2 SAWTOOTH a_13995_11762# VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=700000u
X1371 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1372 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1373 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1374 a_67094_29669# VSS sky130_fd_pr__cap_mim_m3_2 l=1.4e+07u w=1.4e+07u
X1375 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1376 a_11368_10743# a_11080_22588# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1377 a_16885_14913# VREF a_16326_14920# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=900000u
X1378 IL a_11368_10743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1379 a_7812_5796# a_7470_7022# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1380 a_9074_5311# a_7812_5796# a_8654_5311# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X1381 a_81183_36165# a_73231_27552# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X1382 a_71259_32538# a_70429_33459# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X1383 a_7566_10753# a_7278_22598# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1384 VDD IBIAS1 a_16088_14920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1385 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1386 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1387 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1388 VDD IBIAS1 a_16885_14913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=900000u
X1389 a_11168_5307# a_10334_5311# a_10748_5307# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X1390 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1391 a_72247_29498# a_71243_29914# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1392 a_72411_27552# a_56275_30688# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1393 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1394 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1395 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1396 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1397 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1398 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1399 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1400 a_9468_7770# a_8208_7760# a_9048_7770# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=430000u l=150000u
X1401 a_7470_7022# a_14165_10612# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=7.25e+11p pd=5.58e+06u as=0p ps=0u w=2.5e+06u l=500000u
X1402 a_70429_33459# a_66185_27020# a_70439_31826# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1403 VSS a_11368_10743# IL VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1404 VDD a_7566_10753# IL VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1405 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1406 VSS a_66165_10655# a_66125_10752# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1407 a_73011_16066# a_72181_15537# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1408 a_82702_36308# a_82654_36220# OUT VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1409 a_70409_28711# a_69506_31063# a_70419_27078# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1410 IL a_7566_10753# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X1411 a_72177_14863# a_71179_11522# a_72187_13230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
.ends

